package FONT_DEFINITION;

localparam FONT_HEIGHT = 15;
localparam FONT_WIDTH = 8;

/*
localparam logic [0:7] FONT_char0 [0:7] = '{8'h00, 8'hA0, 8'h10, 8'h80, 8'h10, 8'h80, 8'h50, 8'h00};
localparam logic [0:7] FONT_space [0:7] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_exclam [0:7] = '{8'h00, 8'h20, 8'h20, 8'h20, 8'h20, 8'h00, 8'h20, 8'h00};
localparam logic [0:7] FONT_quotedbl [0:7] = '{8'h00, 8'h50, 8'h50, 8'h50, 8'h00, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_numbersign [0:7] = '{8'h50, 8'h50, 8'hF8, 8'h50, 8'hF8, 8'h50, 8'h50, 8'h00};
localparam logic [0:7] FONT_dollar [0:7] = '{8'h20, 8'h70, 8'hA0, 8'h70, 8'h28, 8'h70, 8'h20, 8'h00};
localparam logic [0:7] FONT_percent [0:7] = '{8'h00, 8'h40, 8'h50, 8'h20, 8'h50, 8'h10, 8'h00, 8'h00};
localparam logic [0:7] FONT_ampersand [0:7] = '{8'h40, 8'hA0, 8'hA0, 8'h40, 8'hA0, 8'hA0, 8'h50, 8'h00};
localparam logic [0:7] FONT_quotesingle [0:7] = '{8'h00, 8'h20, 8'h20, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_parenleft [0:7] = '{8'h00, 8'h20, 8'h40, 8'h40, 8'h40, 8'h40, 8'h20, 8'h00};
localparam logic [0:7] FONT_parenright [0:7] = '{8'h00, 8'h40, 8'h20, 8'h20, 8'h20, 8'h20, 8'h40, 8'h00};
localparam logic [0:7] FONT_asterisk [0:7] = '{8'h00, 8'h00, 8'h90, 8'h60, 8'hF0, 8'h60, 8'h90, 8'h00};
localparam logic [0:7] FONT_plus [0:7] = '{8'h00, 8'h00, 8'h20, 8'h20, 8'hF8, 8'h20, 8'h20, 8'h00};
localparam logic [0:7] FONT_comma [0:7] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h30, 8'h20, 8'h40};
localparam logic [0:7] FONT_hyphen [0:7] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'hF0, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_period [0:7] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h70, 8'h20};
localparam logic [0:7] FONT_slash [0:7] = '{8'h00, 8'h10, 8'h10, 8'h20, 8'h40, 8'h80, 8'h80, 8'h00};
localparam logic [0:7] FONT_zero [0:7] = '{8'h00, 8'h20, 8'h50, 8'h50, 8'h50, 8'h50, 8'h20, 8'h00};
localparam logic [0:7] FONT_one [0:7] = '{8'h00, 8'h20, 8'h60, 8'h20, 8'h20, 8'h20, 8'h70, 8'h00};
localparam logic [0:7] FONT_two [0:7] = '{8'h00, 8'h60, 8'h90, 8'h10, 8'h60, 8'h80, 8'hF0, 8'h00};
localparam logic [0:7] FONT_three [0:7] = '{8'h00, 8'hF0, 8'h20, 8'h60, 8'h10, 8'h90, 8'h60, 8'h00};
localparam logic [0:7] FONT_four [0:7] = '{8'h00, 8'h20, 8'h60, 8'hA0, 8'hF0, 8'h20, 8'h20, 8'h00};
localparam logic [0:7] FONT_five [0:7] = '{8'h00, 8'hF0, 8'h80, 8'hE0, 8'h10, 8'h90, 8'h60, 8'h00};
localparam logic [0:7] FONT_six [0:7] = '{8'h00, 8'h60, 8'h80, 8'hE0, 8'h90, 8'h90, 8'h60, 8'h00};
localparam logic [0:7] FONT_seven [0:7] = '{8'h00, 8'hF0, 8'h10, 8'h20, 8'h20, 8'h40, 8'h40, 8'h00};
localparam logic [0:7] FONT_eight [0:7] = '{8'h00, 8'h60, 8'h90, 8'h60, 8'h90, 8'h90, 8'h60, 8'h00};
localparam logic [0:7] FONT_nine [0:7] = '{8'h00, 8'h60, 8'h90, 8'h90, 8'h70, 8'h10, 8'h60, 8'h00};
localparam logic [0:7] FONT_colon [0:7] = '{8'h00, 8'h00, 8'h60, 8'h60, 8'h00, 8'h60, 8'h60, 8'h00};
localparam logic [0:7] FONT_semicolon [0:7] = '{8'h00, 8'h00, 8'h30, 8'h30, 8'h00, 8'h30, 8'h20, 8'h40};
localparam logic [0:7] FONT_less [0:7] = '{8'h00, 8'h10, 8'h20, 8'h40, 8'h40, 8'h20, 8'h10, 8'h00};
localparam logic [0:7] FONT_equal [0:7] = '{8'h00, 8'h00, 8'h00, 8'hF0, 8'h00, 8'hF0, 8'h00, 8'h00};
localparam logic [0:7] FONT_greater [0:7] = '{8'h00, 8'h40, 8'h20, 8'h10, 8'h10, 8'h20, 8'h40, 8'h00};
localparam logic [0:7] FONT_question [0:7] = '{8'h00, 8'h20, 8'h50, 8'h10, 8'h20, 8'h00, 8'h20, 8'h00};
localparam logic [0:7] FONT_at [0:7] = '{8'h30, 8'h48, 8'h98, 8'hA8, 8'hA8, 8'h90, 8'h40, 8'h30};
localparam logic [0:7] FONT_A [0:7] = '{8'h00, 8'h60, 8'h90, 8'h90, 8'hF0, 8'h90, 8'h90, 8'h00};
localparam logic [0:7] FONT_B [0:7] = '{8'h00, 8'hE0, 8'h90, 8'hE0, 8'h90, 8'h90, 8'hE0, 8'h00};
localparam logic [0:7] FONT_C [0:7] = '{8'h00, 8'h60, 8'h90, 8'h80, 8'h80, 8'h90, 8'h60, 8'h00};
localparam logic [0:7] FONT_D [0:7] = '{8'h00, 8'hE0, 8'h90, 8'h90, 8'h90, 8'h90, 8'hE0, 8'h00};
localparam logic [0:7] FONT_E [0:7] = '{8'h00, 8'hF0, 8'h80, 8'hE0, 8'h80, 8'h80, 8'hF0, 8'h00};
localparam logic [0:7] FONT_F [0:7] = '{8'h00, 8'hF0, 8'h80, 8'hE0, 8'h80, 8'h80, 8'h80, 8'h00};
localparam logic [0:7] FONT_G [0:7] = '{8'h00, 8'h60, 8'h90, 8'h80, 8'hB0, 8'h90, 8'h60, 8'h00};
localparam logic [0:7] FONT_H [0:7] = '{8'h00, 8'h90, 8'h90, 8'hF0, 8'h90, 8'h90, 8'h90, 8'h00};
localparam logic [0:7] FONT_I [0:7] = '{8'h00, 8'h70, 8'h20, 8'h20, 8'h20, 8'h20, 8'h70, 8'h00};
localparam logic [0:7] FONT_J [0:7] = '{8'h00, 8'h70, 8'h20, 8'h20, 8'h20, 8'hA0, 8'h40, 8'h00};
localparam logic [0:7] FONT_K [0:7] = '{8'h00, 8'h90, 8'hA0, 8'hC0, 8'hA0, 8'hA0, 8'h90, 8'h00};
localparam logic [0:7] FONT_L [0:7] = '{8'h00, 8'h80, 8'h80, 8'h80, 8'h80, 8'h80, 8'hF0, 8'h00};
localparam logic [0:7] FONT_M [0:7] = '{8'h00, 8'h90, 8'hF0, 8'hF0, 8'h90, 8'h90, 8'h90, 8'h00};
localparam logic [0:7] FONT_N [0:7] = '{8'h00, 8'h90, 8'hD0, 8'hF0, 8'hB0, 8'hB0, 8'h90, 8'h00};
localparam logic [0:7] FONT_O [0:7] = '{8'h00, 8'h60, 8'h90, 8'h90, 8'h90, 8'h90, 8'h60, 8'h00};
localparam logic [0:7] FONT_P [0:7] = '{8'h00, 8'hE0, 8'h90, 8'h90, 8'hE0, 8'h80, 8'h80, 8'h00};
localparam logic [0:7] FONT_Q [0:7] = '{8'h00, 8'h60, 8'h90, 8'h90, 8'hD0, 8'hB0, 8'h60, 8'h10};
localparam logic [0:7] FONT_R [0:7] = '{8'h00, 8'hE0, 8'h90, 8'h90, 8'hE0, 8'h90, 8'h90, 8'h00};
localparam logic [0:7] FONT_S [0:7] = '{8'h00, 8'h60, 8'h90, 8'h40, 8'h20, 8'h90, 8'h60, 8'h00};
localparam logic [0:7] FONT_T [0:7] = '{8'h00, 8'h70, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h00};
localparam logic [0:7] FONT_U [0:7] = '{8'h00, 8'h90, 8'h90, 8'h90, 8'h90, 8'h90, 8'h60, 8'h00};
localparam logic [0:7] FONT_V [0:7] = '{8'h00, 8'h90, 8'h90, 8'h90, 8'h90, 8'h60, 8'h60, 8'h00};
localparam logic [0:7] FONT_W [0:7] = '{8'h00, 8'h90, 8'h90, 8'h90, 8'hF0, 8'hF0, 8'h90, 8'h00};
localparam logic [0:7] FONT_X [0:7] = '{8'h00, 8'h90, 8'h90, 8'h60, 8'h60, 8'h90, 8'h90, 8'h00};
localparam logic [0:7] FONT_Y [0:7] = '{8'h00, 8'h88, 8'h88, 8'h50, 8'h20, 8'h20, 8'h20, 8'h00};
localparam logic [0:7] FONT_Z [0:7] = '{8'h00, 8'hF0, 8'h10, 8'h20, 8'h40, 8'h80, 8'hF0, 8'h00};
localparam logic [0:7] FONT_bracketleft [0:7] = '{8'h00, 8'h70, 8'h40, 8'h40, 8'h40, 8'h40, 8'h70, 8'h00};
localparam logic [0:7] FONT_backslash [0:7] = '{8'h00, 8'h80, 8'h80, 8'h40, 8'h20, 8'h10, 8'h10, 8'h00};
localparam logic [0:7] FONT_bracketright [0:7] = '{8'h00, 8'h70, 8'h10, 8'h10, 8'h10, 8'h10, 8'h70, 8'h00};
localparam logic [0:7] FONT_asciicircum [0:7] = '{8'h00, 8'h20, 8'h50, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_underscore [0:7] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hF0};
localparam logic [0:7] FONT_grave [0:7] = '{8'h00, 8'h40, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_a [0:7] = '{8'h00, 8'h00, 8'h00, 8'h70, 8'h90, 8'h90, 8'h70, 8'h00};
localparam logic [0:7] FONT_b [0:7] = '{8'h00, 8'h80, 8'h80, 8'hE0, 8'h90, 8'h90, 8'hE0, 8'h00};
localparam logic [0:7] FONT_c [0:7] = '{8'h00, 8'h00, 8'h00, 8'h30, 8'h40, 8'h40, 8'h30, 8'h00};
localparam logic [0:7] FONT_d [0:7] = '{8'h00, 8'h10, 8'h10, 8'h70, 8'h90, 8'h90, 8'h70, 8'h00};
localparam logic [0:7] FONT_e [0:7] = '{8'h00, 8'h00, 8'h00, 8'h60, 8'hB0, 8'hC0, 8'h60, 8'h00};
localparam logic [0:7] FONT_f [0:7] = '{8'h00, 8'h20, 8'h50, 8'h40, 8'hE0, 8'h40, 8'h40, 8'h00};
localparam logic [0:7] FONT_g [0:7] = '{8'h00, 8'h00, 8'h00, 8'h60, 8'h90, 8'h70, 8'h10, 8'h60};
localparam logic [0:7] FONT_h [0:7] = '{8'h00, 8'h80, 8'h80, 8'hE0, 8'h90, 8'h90, 8'h90, 8'h00};
localparam logic [0:7] FONT_i [0:7] = '{8'h00, 8'h20, 8'h00, 8'h60, 8'h20, 8'h20, 8'h70, 8'h00};
localparam logic [0:7] FONT_j [0:7] = '{8'h00, 8'h10, 8'h00, 8'h10, 8'h10, 8'h10, 8'h50, 8'h20};
localparam logic [0:7] FONT_k [0:7] = '{8'h00, 8'h80, 8'h80, 8'h90, 8'hE0, 8'h90, 8'h90, 8'h00};
localparam logic [0:7] FONT_l [0:7] = '{8'h00, 8'h60, 8'h20, 8'h20, 8'h20, 8'h20, 8'h70, 8'h00};
localparam logic [0:7] FONT_m [0:7] = '{8'h00, 8'h00, 8'h00, 8'hD0, 8'hA8, 8'hA8, 8'hA8, 8'h00};
localparam logic [0:7] FONT_n [0:7] = '{8'h00, 8'h00, 8'h00, 8'hE0, 8'h90, 8'h90, 8'h90, 8'h00};
localparam logic [0:7] FONT_o [0:7] = '{8'h00, 8'h00, 8'h00, 8'h60, 8'h90, 8'h90, 8'h60, 8'h00};
localparam logic [0:7] FONT_p [0:7] = '{8'h00, 8'h00, 8'h00, 8'hE0, 8'h90, 8'hE0, 8'h80, 8'h80};
localparam logic [0:7] FONT_q [0:7] = '{8'h00, 8'h00, 8'h00, 8'h70, 8'h90, 8'h70, 8'h10, 8'h10};
localparam logic [0:7] FONT_r [0:7] = '{8'h00, 8'h00, 8'h00, 8'hA0, 8'hD0, 8'h80, 8'h80, 8'h00};
localparam logic [0:7] FONT_s [0:7] = '{8'h00, 8'h00, 8'h00, 8'h30, 8'h60, 8'h10, 8'h60, 8'h00};
localparam logic [0:7] FONT_t [0:7] = '{8'h00, 8'h40, 8'h40, 8'hE0, 8'h40, 8'h50, 8'h20, 8'h00};
localparam logic [0:7] FONT_u [0:7] = '{8'h00, 8'h00, 8'h00, 8'h90, 8'h90, 8'h90, 8'h70, 8'h00};
localparam logic [0:7] FONT_v [0:7] = '{8'h00, 8'h00, 8'h00, 8'h50, 8'h50, 8'h50, 8'h20, 8'h00};
localparam logic [0:7] FONT_w [0:7] = '{8'h00, 8'h00, 8'h00, 8'h88, 8'hA8, 8'hA8, 8'h50, 8'h00};
localparam logic [0:7] FONT_x [0:7] = '{8'h00, 8'h00, 8'h00, 8'h90, 8'h60, 8'h60, 8'h90, 8'h00};
localparam logic [0:7] FONT_y [0:7] = '{8'h00, 8'h00, 8'h00, 8'h90, 8'h90, 8'h70, 8'h90, 8'h60};
localparam logic [0:7] FONT_z [0:7] = '{8'h00, 8'h00, 8'h00, 8'hF0, 8'h20, 8'h40, 8'hF0, 8'h00};
*/

localparam logic [0:7] FONT_char0 [0:14] = '{8'h00, 8'h00, 8'h6D, 8'h01, 8'h40, 8'h41, 8'h01, 8'h40, 8'h41, 8'h01, 8'h40, 8'h5B, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_space [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_exclam [0:14] = '{8'h00, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h00, 8'h00, 8'h08, 8'h08, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_quotedbl [0:14] = '{8'h00, 8'h00, 8'h12, 8'h12, 8'h12, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_numbersign [0:14] = '{8'h00, 8'h00, 8'h00, 8'h24, 8'h24, 8'h7E, 8'h24, 8'h24, 8'h7E, 8'h24, 8'h24, 8'h00, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_dollar [0:14] = '{8'h00, 8'h00, 8'h08, 8'h3E, 8'h49, 8'h48, 8'h28, 8'h1C, 8'h0A, 8'h09, 8'h49, 8'h3E, 8'h08, 8'h00, 8'h00};
localparam logic [0:7] FONT_percent [0:14] = '{8'h00, 8'h00, 8'h21, 8'h52, 8'h52, 8'h24, 8'h08, 8'h08, 8'h12, 8'h25, 8'h25, 8'h42, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_ampersand [0:14] = '{8'h00, 8'h00, 8'h30, 8'h48, 8'h48, 8'h48, 8'h30, 8'h31, 8'h4A, 8'h44, 8'h4A, 8'h31, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_quotesingle [0:14] = '{8'h00, 8'h00, 8'h08, 8'h08, 8'h08, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_parenleft [0:14] = '{8'h00, 8'h04, 8'h08, 8'h08, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h08, 8'h08, 8'h04, 8'h00, 8'h00};
localparam logic [0:7] FONT_parenright [0:14] = '{8'h00, 8'h10, 8'h08, 8'h08, 8'h04, 8'h04, 8'h04, 8'h04, 8'h04, 8'h04, 8'h08, 8'h08, 8'h10, 8'h00, 8'h00};
localparam logic [0:7] FONT_asterisk [0:14] = '{8'h00, 8'h00, 8'h08, 8'h49, 8'h2A, 8'h1C, 8'h2A, 8'h49, 8'h08, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_plus [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h08, 8'h08, 8'h08, 8'h7F, 8'h08, 8'h08, 8'h08, 8'h00, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_comma [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0C, 8'h0C, 8'h04, 8'h04, 8'h08};
localparam logic [0:7] FONT_hyphen [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_period [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0C, 8'h0C, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_slash [0:14] = '{8'h00, 8'h00, 8'h01, 8'h02, 8'h02, 8'h04, 8'h08, 8'h08, 8'h10, 8'h20, 8'h20, 8'h40, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_zero [0:14] = '{8'h00, 8'h00, 8'h1C, 8'h22, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h22, 8'h1C, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_one [0:14] = '{8'h00, 8'h00, 8'h08, 8'h18, 8'h28, 8'h48, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h7F, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_two [0:14] = '{8'h00, 8'h00, 8'h3E, 8'h41, 8'h41, 8'h02, 8'h04, 8'h08, 8'h10, 8'h20, 8'h40, 8'h7F, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_three [0:14] = '{8'h00, 8'h00, 8'h7F, 8'h01, 8'h02, 8'h04, 8'h0E, 8'h01, 8'h01, 8'h01, 8'h41, 8'h3E, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_four [0:14] = '{8'h00, 8'h00, 8'h02, 8'h06, 8'h0A, 8'h12, 8'h22, 8'h42, 8'h7F, 8'h02, 8'h02, 8'h02, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_five [0:14] = '{8'h00, 8'h00, 8'h7F, 8'h40, 8'h40, 8'h5E, 8'h61, 8'h01, 8'h01, 8'h01, 8'h41, 8'h3E, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_six [0:14] = '{8'h00, 8'h00, 8'h1E, 8'h20, 8'h40, 8'h40, 8'h5E, 8'h61, 8'h41, 8'h41, 8'h41, 8'h3E, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_seven [0:14] = '{8'h00, 8'h00, 8'h7F, 8'h01, 8'h02, 8'h02, 8'h04, 8'h04, 8'h08, 8'h08, 8'h10, 8'h10, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_eight [0:14] = '{8'h00, 8'h00, 8'h1C, 8'h22, 8'h41, 8'h22, 8'h1C, 8'h22, 8'h41, 8'h41, 8'h22, 8'h1C, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_nine [0:14] = '{8'h00, 8'h00, 8'h3E, 8'h41, 8'h41, 8'h41, 8'h43, 8'h3D, 8'h01, 8'h01, 8'h02, 8'h3C, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_colon [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0C, 8'h0C, 8'h00, 8'h00, 8'h00, 8'h0C, 8'h0C, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_semicolon [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h0C, 8'h0C, 8'h00, 8'h00, 8'h00, 8'h0C, 8'h0C, 8'h04, 8'h04, 8'h08};
localparam logic [0:7] FONT_less [0:14] = '{8'h00, 8'h00, 8'h02, 8'h04, 8'h08, 8'h10, 8'h20, 8'h20, 8'h10, 8'h08, 8'h04, 8'h02, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_equal [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7F, 8'h00, 8'h00, 8'h7F, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_greater [0:14] = '{8'h00, 8'h00, 8'h20, 8'h10, 8'h08, 8'h04, 8'h02, 8'h02, 8'h04, 8'h08, 8'h10, 8'h20, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_question [0:14] = '{8'h00, 8'h00, 8'h3E, 8'h41, 8'h41, 8'h01, 8'h02, 8'h04, 8'h08, 8'h08, 8'h00, 8'h08, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_at [0:14] = '{8'h00, 8'h00, 8'h3E, 8'h41, 8'h41, 8'h4F, 8'h51, 8'h53, 8'h4D, 8'h40, 8'h40, 8'h3E, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_A [0:14] = '{8'h00, 8'h00, 8'h08, 8'h14, 8'h22, 8'h41, 8'h41, 8'h41, 8'h7F, 8'h41, 8'h41, 8'h41, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_B [0:14] = '{8'h00, 8'h00, 8'h7C, 8'h42, 8'h41, 8'h42, 8'h7C, 8'h42, 8'h41, 8'h41, 8'h42, 8'h7C, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_C [0:14] = '{8'h00, 8'h00, 8'h3E, 8'h41, 8'h40, 8'h40, 8'h40, 8'h40, 8'h40, 8'h40, 8'h41, 8'h3E, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_D [0:14] = '{8'h00, 8'h00, 8'h7C, 8'h42, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h42, 8'h7C, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_E [0:14] = '{8'h00, 8'h00, 8'h7F, 8'h40, 8'h40, 8'h40, 8'h7C, 8'h40, 8'h40, 8'h40, 8'h40, 8'h7F, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_F [0:14] = '{8'h00, 8'h00, 8'h7F, 8'h40, 8'h40, 8'h40, 8'h7C, 8'h40, 8'h40, 8'h40, 8'h40, 8'h40, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_G [0:14] = '{8'h00, 8'h00, 8'h3E, 8'h41, 8'h40, 8'h40, 8'h40, 8'h47, 8'h41, 8'h41, 8'h41, 8'h3E, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_H [0:14] = '{8'h00, 8'h00, 8'h41, 8'h41, 8'h41, 8'h41, 8'h7F, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_I [0:14] = '{8'h00, 8'h00, 8'h3E, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h3E, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_J [0:14] = '{8'h00, 8'h00, 8'h0F, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02, 8'h42, 8'h3C, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_K [0:14] = '{8'h00, 8'h00, 8'h41, 8'h42, 8'h44, 8'h48, 8'h70, 8'h50, 8'h48, 8'h44, 8'h42, 8'h41, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_L [0:14] = '{8'h00, 8'h00, 8'h40, 8'h40, 8'h40, 8'h40, 8'h40, 8'h40, 8'h40, 8'h40, 8'h40, 8'h7F, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_M [0:14] = '{8'h00, 8'h00, 8'h41, 8'h41, 8'h63, 8'h55, 8'h55, 8'h49, 8'h49, 8'h41, 8'h41, 8'h41, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_N [0:14] = '{8'h00, 8'h00, 8'h41, 8'h41, 8'h61, 8'h51, 8'h49, 8'h45, 8'h43, 8'h41, 8'h41, 8'h41, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_O [0:14] = '{8'h00, 8'h00, 8'h3E, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h3E, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_P [0:14] = '{8'h00, 8'h00, 8'h7E, 8'h41, 8'h41, 8'h41, 8'h7E, 8'h40, 8'h40, 8'h40, 8'h40, 8'h40, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_Q [0:14] = '{8'h00, 8'h00, 8'h3E, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h51, 8'h49, 8'h3E, 8'h04, 8'h03, 8'h00};
localparam logic [0:7] FONT_R [0:14] = '{8'h00, 8'h00, 8'h7E, 8'h41, 8'h41, 8'h41, 8'h7E, 8'h48, 8'h44, 8'h42, 8'h41, 8'h41, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_S [0:14] = '{8'h00, 8'h00, 8'h3E, 8'h41, 8'h41, 8'h40, 8'h38, 8'h06, 8'h01, 8'h41, 8'h41, 8'h3E, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_T [0:14] = '{8'h00, 8'h00, 8'h7F, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_U [0:14] = '{8'h00, 8'h00, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h3E, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_V [0:14] = '{8'h00, 8'h00, 8'h41, 8'h41, 8'h41, 8'h22, 8'h22, 8'h22, 8'h14, 8'h14, 8'h14, 8'h08, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_W [0:14] = '{8'h00, 8'h00, 8'h41, 8'h41, 8'h41, 8'h41, 8'h49, 8'h49, 8'h49, 8'h49, 8'h55, 8'h22, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_X [0:14] = '{8'h00, 8'h00, 8'h41, 8'h41, 8'h22, 8'h14, 8'h08, 8'h08, 8'h14, 8'h22, 8'h41, 8'h41, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_Y [0:14] = '{8'h00, 8'h00, 8'h41, 8'h41, 8'h22, 8'h14, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_Z [0:14] = '{8'h00, 8'h00, 8'h7F, 8'h01, 8'h02, 8'h04, 8'h08, 8'h10, 8'h20, 8'h40, 8'h40, 8'h7F, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_bracketleft [0:14] = '{8'h00, 8'h1E, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h10, 8'h1E, 8'h00, 8'h00};
localparam logic [0:7] FONT_backslash [0:14] = '{8'h00, 8'h00, 8'h40, 8'h20, 8'h20, 8'h10, 8'h08, 8'h08, 8'h04, 8'h02, 8'h02, 8'h01, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_bracketright [0:14] = '{8'h00, 8'h3C, 8'h04, 8'h04, 8'h04, 8'h04, 8'h04, 8'h04, 8'h04, 8'h04, 8'h04, 8'h04, 8'h3C, 8'h00, 8'h00};
localparam logic [0:7] FONT_asciicircum [0:14] = '{8'h00, 8'h00, 8'h08, 8'h14, 8'h22, 8'h41, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_underscore [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h00};
localparam logic [0:7] FONT_grave [0:14] = '{8'h00, 8'h10, 8'h08, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_a [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3E, 8'h01, 8'h01, 8'h3F, 8'h41, 8'h43, 8'h3D, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_b [0:14] = '{8'h00, 8'h00, 8'h40, 8'h40, 8'h40, 8'h5E, 8'h61, 8'h41, 8'h41, 8'h41, 8'h61, 8'h5E, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_c [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3E, 8'h41, 8'h40, 8'h40, 8'h40, 8'h41, 8'h3E, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_d [0:14] = '{8'h00, 8'h00, 8'h01, 8'h01, 8'h01, 8'h3D, 8'h43, 8'h41, 8'h41, 8'h41, 8'h43, 8'h3D, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_e [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3E, 8'h41, 8'h41, 8'h7F, 8'h40, 8'h40, 8'h3E, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_f [0:14] = '{8'h00, 8'h00, 8'h0E, 8'h11, 8'h11, 8'h10, 8'h10, 8'h7C, 8'h10, 8'h10, 8'h10, 8'h10, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_g [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3D, 8'h42, 8'h42, 8'h42, 8'h3C, 8'h40, 8'h3E, 8'h41, 8'h41, 8'h3E};
localparam logic [0:7] FONT_h [0:14] = '{8'h00, 8'h00, 8'h40, 8'h40, 8'h40, 8'h5E, 8'h61, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_i [0:14] = '{8'h00, 8'h00, 8'h18, 8'h00, 8'h00, 8'h38, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h3E, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_j [0:14] = '{8'h00, 8'h00, 8'h06, 8'h00, 8'h00, 8'h0E, 8'h02, 8'h02, 8'h02, 8'h02, 8'h02, 8'h42, 8'h42, 8'h42, 8'h3C};
localparam logic [0:7] FONT_k [0:14] = '{8'h00, 8'h00, 8'h40, 8'h40, 8'h40, 8'h41, 8'h46, 8'h58, 8'h60, 8'h58, 8'h46, 8'h41, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_l [0:14] = '{8'h00, 8'h00, 8'h38, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h08, 8'h3E, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_m [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h76, 8'h49, 8'h49, 8'h49, 8'h49, 8'h49, 8'h41, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_n [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h5E, 8'h61, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_o [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3E, 8'h41, 8'h41, 8'h41, 8'h41, 8'h41, 8'h3E, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_p [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h5E, 8'h61, 8'h41, 8'h41, 8'h41, 8'h61, 8'h5E, 8'h40, 8'h40, 8'h40};
localparam logic [0:7] FONT_q [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3D, 8'h43, 8'h41, 8'h41, 8'h41, 8'h43, 8'h3D, 8'h01, 8'h01, 8'h01};
localparam logic [0:7] FONT_r [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h4E, 8'h31, 8'h21, 8'h20, 8'h20, 8'h20, 8'h20, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_s [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h3E, 8'h41, 8'h40, 8'h3E, 8'h01, 8'h41, 8'h3E, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_t [0:14] = '{8'h00, 8'h00, 8'h00, 8'h10, 8'h10, 8'h7E, 8'h10, 8'h10, 8'h10, 8'h10, 8'h11, 8'h0E, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_u [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h42, 8'h42, 8'h42, 8'h42, 8'h42, 8'h42, 8'h3D, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_v [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h41, 8'h41, 8'h22, 8'h22, 8'h14, 8'h14, 8'h08, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_w [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h41, 8'h41, 8'h49, 8'h49, 8'h49, 8'h55, 8'h22, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_x [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h41, 8'h22, 8'h14, 8'h08, 8'h14, 8'h22, 8'h41, 8'h00, 8'h00, 8'h00};
localparam logic [0:7] FONT_y [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h42, 8'h42, 8'h42, 8'h42, 8'h42, 8'h46, 8'h3A, 8'h02, 8'h42, 8'h3C};
localparam logic [0:7] FONT_z [0:14] = '{8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h7F, 8'h02, 8'h04, 8'h08, 8'h10, 8'h20, 8'h7F, 8'h00, 8'h00, 8'h00};

endpackage
