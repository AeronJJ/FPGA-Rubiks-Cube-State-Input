`timescale 1ns / 100ps
module TEXT_GENERATOR_tb;

reg en = 1'b1;
reg [8:0] x_pixel = 9'b0;
reg [7:0] y_pixel = 8'b0;
wire [15:0] pixel;
wire active;

TEXT_GENERATOR #(.size(1)) dut (
	en,
	x_pixel,
	y_pixel,
	pixel,
	active
);

always #5 begin
	if (y_pixel == 8'd240) begin
		y_pixel <= 1'b0;
		x_pixel <= 1'b0;
	end
	else if (x_pixel == 9'd320) begin
		x_pixel <= 1'b0;
		y_pixel <= y_pixel + 1'b1;
	end
	else begin
		x_pixel <= x_pixel + 1'b1;
	end
end

//initial begin
	
//end

endmodule
