package MSP2807_COLOURS;

localparam MSP_WHITE 	= 16'hFFFF;
localparam MSP_BLACK 	= 16'h0000;
localparam MSP_RED 		= 16'hF800;
localparam MSP_BLUE 		= 16'h001F;
localparam MSP_GREEN 	= 16'h07E0;
localparam MSP_ORANGE 	= 16'hFD68;
localparam MSP_YELLOW 	= 16'hFFC0;

endpackage
